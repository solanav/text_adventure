#o:1|Torch|-1|Lights your way|1|0|-1|1|0|
#o:2|Key1|13|Just a broken fragment|1|0|-1|0|0|
#o:3|Key2|53|Just a broken fragment|1|0|-1|0|0|
#o:4|Key3|65|Just a broken fragment|1|0|-1|0|0|
#o:5|Key4|26|Just a broken fragment|1|0|-1|0|0|
#o:6|Key5|45|Just a broken fragment|1|0|-1|0|0|
#o:7|Note1|13|Note 1 description|0|0|-1|0|0|
#o:8|Note2|53|Note 2 description|0|0|-1|0|0|
#o:9|Note3|65|Note 3 description|0|0|-1|0|0|
#o:10|Note4|26|Note 4 description|0|0|-1|0|0|
#o:11|Note5|45|Note 5 description|0|0|-1|0|0|
#o:12|Bottle|25|There's a sticky substance|1|0|-1|0|0|
#o:13|RockXL|66|It's got big bones|0|0|0|0|0|
#o:14|RockM|15|Do you know big rock?|0|0|0|0|0|
#o:15|RockS|11|Do you know medium rock?|0|0|0|0|0|
#o:16|Stick|25|Why would you take it?|0|0|0|0|0|
#o:17|Leafs|-1||0|0|0|0|0|
#o:18|Tree|35|Yeah, a tree|0|0|0|0|0|
#o:19|Wand|42|You are no wizard Dante!|0|0|-1|0|0|
#o:20|Sword|42|You are no warrior Dante!|0|0|-1|0|0|
#o:21|MasterKey|16|That wasn't that hard was it?|1|0|62|0|0|
#p:1|
#l:1|Link 1|11|12|0|0|
#l:2|Link 2|12|11|2|0|
#l:3|Link 3|12|13|0|0|
#l:4|Link 4|13|12|2|0|
#l:5|Link 5|13|14|0|0|
#l:6|Link 6|14|13|2|0|
#l:7|Link 7|14|15|0|0|
#l:8|Link 8|15|14|2|0|
#l:9|Link 9|21|22|0|0|
#l:10|Link 10|22|21|2|0|
#l:11|Link 11|22|23|0|0|
#l:12|Link 12|23|22|2|0|
#l:13|Link 13|23|24|0|0|
#l:14|Link 14|24|23|2|0|
#l:15|Link 15|24|25|0|0|
#l:16|Link 16|25|24|2|0|
#l:17|Link 17|25|26|0|0|
#l:18|Link 18|26|25|2|0|
#l:19|Link 19|41|42|0|0|
#l:20|Link 20|42|41|2|0|
#l:21|Link 21|42|43|0|0|
#l:22|Link 22|43|42|2|0|
#l:23|Link 23|51|52|0|0|
#l:24|Link 24|52|51|2|0|
#l:25|Link 25|52|53|0|0|
#l:26|Link 26|53|52|2|0|
#l:27|Link 27|53|54|0|0|
#l:28|Link 28|54|53|2|0|
#l:29|Link 29|54|55|0|0|
#l:30|Link 30|55|54|2|0|
#l:31|Link 31|55|56|0|0|
#l:32|Link 32|56|55|2|0|
#l:33|Link 33|64|65|0|0|
#l:34|Link 34|65|64|2|0|
#l:35|Link 35|65|66|0|0|
#l:36|Link 36|66|65|2|0|
#l:37|Link 37|11|21|1|0|
#l:38|Link 38|21|11|3|0|
#l:39|Link 39|21|31|1|0|
#l:40|Link 40|31|21|3|0|
#l:41|Link 41|31|41|1|0|
#l:42|Link 42|41|31|3|0|
#l:43|Link 43|41|51|1|0|
#l:44|Link 44|51|41|3|0|
#l:45|Link 45|52|62|1|0|
#l:46|Link 46|62|52|3|0|
#l:47|Link 47|23|33|1|0|
#l:48|Link 48|33|23|3|0|
#l:49|Link 49|33|43|1|0|
#l:50|Link 50|43|33|3|0|
#l:51|Link 51|44|54|1|0|
#l:52|Link 52|54|44|3|0|
#l:53|Link 53|54|64|1|0|
#l:54|Link 54|64|54|3|0|
#l:55|Link 55|15|25|1|0|
#l:56|Link 56|25|15|3|0|
#l:57|Link 57|25|35|1|0|
#l:58|Link 58|35|25|3|0|
#l:59|Link 59|35|45|1|0|
#l:60|Link 60|45|35|3|0|
#l:61|Link 61|26|36|1|0|
#l:62|Link 62|36|26|3|0|
#l:63|Link 63|36|46|1|0|
#l:64|Link 64|46|36|3|0|
#l:65|Link 65|46|56|1|0|
#l:66|Link 66|56|46|3|0|
#l:67|Link 67|56|66|1|0|
#l:68|Link 68|66|56|3|0|
#l:69|Link 69|35|36|0|0|
#l:70|Link 70|36|35|2|0|
#l:71|Link 71|36|25|0|0|
#l:72|Link 72|44|45|0|0|
#l:73|Link 73|45|44|2|0|
#l:74|Link 74|62|61|2|1|
