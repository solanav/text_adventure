�D            ��E    saves/hay.sv    
       �w@     ����   H�            �    �w@     ���            ����   ����    ���u�У@���   �j@     `���   �D     hay    �D       	         save                            hay                             save hay ���u�У`���   a@     �D     �D      ���   �@     ����   ���           �D     �D     `�,    hr@     sr@     {r@     �r@     �r@     �r@     �r@     �r@     ./log/                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          �q@      ���u�У����           �q@     0��            ����   �\"   V@             �u���0�`@     ����                   ����$/��e%��0�                       Pr@     �
    �                    �K     ����   `@      ���u�У����   �@     ����   �D            ��E    saves/hay.sv    
       �w@     ����   H�            �    �w@     ���            ����   ����    ���u�У@���   �j@     `���   �D     hay    �D       	         save                            hay                             save hay ���u�У`���   a@     �D     �D      ���   �@     ����   ���           �D     �D     `�,    hr@     sr@     {r@     �r@     �r@     �r@     �r@     �r@     ./log/                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   P     `@        �$     ���u�У����   �@     ����   �D            ��E    saves/hay.sv    
       �w@     ����   H�            �    �w@     ���            ����   ����    ���u�У@���   �j@     `���   �D     hay    �D       	         save                            hay                             save hay ���u�У`���   a@     �D     �D      ���   �@     ����   ���           �D     �D     `�,    hr@     sr@     {r@     �r@     �r@     �r@     �r@     �r@     ./log/                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          �q@      ���u�У����           �q@     0��            ����   �\"   V@             �u���0�`@     ����                   ����$/��e%��0�                       Pr@     �
    �                    `@     ����           �@     ����                 ����   ����           ����   ����   ����     �   '  �   W  �   d  �   n  �   }  �   �  �   �  �   �  �   �  �   �  �   �  �    �   K �   � �   � �   � �    �   > �   r �   � �   � �   � �   ? �   J �   i �   � �   � �   � �   � �      ��     �$     ���u�У����   �@     ����   �D            ��E    saves/hay.sv    
       �w@     ����   H�            �    �w@     ���            ����   ����    ���u�У@���   �j@     `���   �D     hay    �D       	         save                            hay                             save hay ���u�У`���   a@     �D     �D      ���   �@     ����   ���           �D     �D     `�,    hr@     sr@     {r@     �r@     �r@     �r@     �r@     �r@     ./log/                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          �q@      ���u�У����           �q@     0��            ����   �\"   V@             �u���0�`@     ����                   ����$/��e%��0�                       Pr@     �
    �                    `@     ����           �@     ����                 ����   ����           ����   ����   ����     �   '  �   W  �   d  �   n  �   }  �   �  �   �  �   �  �   �  �   �  �   �  �    �   K �   � �   � �   � �    �   > �   r �   � �   � �   � �   ? �   J �   i �   � �   � �   � �   � �   
 �    �   3 �   S �   b �   � �   `�E     ���u�У����   �@     ����   �D            ��E    saves/hay.sv    
       �w@     ����   H�            �    �w@     ���            ����   ����    ���u�У@���   �j@     `���   �D     hay    �D       	         save                            hay                             save hay ���u�У`���   a@     �D     �D      ���   �@     ����   ���           �D     �D     `�,    hr@     sr@     {r@     �r@     �r@     �r@     �r@     �r@     ./log/                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          �q@      ���u�У����           �q@     0��            ����   �\"   V@             �u���0�`@     ����                   ����$/��e%��0�                       Pr@     �
    �                    `@     ����           �@     ����                 ����   ����           ����   ����   ����     �   '  �   W  �   d  �   n  �   }  �   �  �   �  �   �  �   �  �   �  �   �  �    �   K �   � �   � �   � �    �   > �   r �   � �   � �   � �   ? �   J �   i �   � �   � �   � �   � �   
 �    �   3 �   S �   b �   � �   � �   � �     �   � �    �   ; �   O �   n �   � �   � �   � �   � �   � �   � �   � �    �   � �   � �   � �   � �    �   1 �   I �   \ �   ~ �   � �   � �   � �   � �   � �    �   � �    �   ' �   / �   D �   Y �   m �                   0.��         ���                         d              @ @            8              	                                    	       `@            �             �             �             �                            � �          � �          � �                                      ./game_exec data.dat LESSOPEN=| /usr/bin/lesspipe %s PROFILEHOME= KDE_FULL_SESSION=true GS_LIB=/home/krantup/.fonts PAM_KWALLET5_LOGIN=/tmp/kwallet5_krantup.socket USER=krantup LANGUAGE= XDG_SEAT=seat0 XDG_SESSION_TYPE=x11 SSH_AGENT_PID=1309 XCURSOR_SIZE=0 SHLVL=1 LD_LIBRARY_PATH=/usr/lib/debug HOME=/home/krantup OLDPWD=/home/krantup/like_ocas_in_the_rain/saves DESKTOP_SESSION=/usr/share/xsessions/plasma XDG_SESSION_COOKIE=f06880154fba4ddd9dd7dbf4157fe0d9-1523966234.406189-1737042203 GTK_RC_FILES=/etc/gtk/gtkrc:/home/krantup/.gtkrc:/home/krantup/.config/gtkrc KDE_SESSION_VERSION=5 GTK_MODULES=gail:atk-bridge QT_LINUX_ACCESSIBILITY_ALWAYS_ON=1 XDG_SEAT_PATH=/org/freedesktop/DisplayManager/Seat0 SHELL_SESSION_ID=611bf9cdea254000a7042aeb286587d4 KONSOLE_DBUS_SESSION=/Sessions/1 LC_MONETARY=es_ES.UTF-8 DBUS_SESSION_BUS_ADDRESS=unix:abstract=/tmp/dbus-reuyjzkE9j,guid=c717f1e3ead3d5c0396501d75ad5e11a MAKEFLAGS= KONSOLE_DBUS_WINDOW=/Windows/1 MAKE_TERMERR=/dev/pts/1 MANDATORY_PATH=/usr/share/gconf//usr/share/xsessions/plasma.mandatory.path LOGNAME=krantup _=/usr/bin/make QT_AUTO_SCREEN_SCALE_FACTOR=0 WINDOWID=10485765 XDG_SESSION_CLASS=user KONSOLE_PROFILE_NAME=Linux Mint COLORFGBG=15;0 DEFAULTS_PATH=/usr/share/gconf//usr/share/xsessions/plasma.default.path XDG_SESSION_ID=2 TERM=xterm GTK2_RC_FILES=/etc/gtk-2.0/gtkrc:/home/krantup/.gtkrc-2.0:/home/krantup/.config/gtkrc-2.0 PATH=/home/krantup/bin:/home/krantup/.local/bin:/usr/local/sbin:/usr/local/bin:/usr/sbin:/usr/bin:/sbin:/bin:/usr/games:/usr/local/games SESSION_MANAGER=local/kde-mint1:@/tmp/.ICE-unix/1638,unix/kde-mint1:/tmp/.ICE-unix/1638 XDG_SESSION_PATH=/org/freedesktop/DisplayManager/Session1 XCURSOR_THEME=Bread XDG_RUNTIME_DIR=/run/user/1000 LC_ADDRESS=es_ES.UTF-8 MAKELEVEL=1 GLIBCPP_FORCE_NEW=1 DISPLAY=:0 XDG_CURRENT_DESKTOP=KDE LC_TELEPHONE=es_ES.UTF-8 LANG=en_US.UTF-8 XAUTHORITY=/tmp/xauth-1000-_0 LS_COLORS=rs=0:di=01;34:ln=01;36:mh=00:pi=40;33:so=01;35:do=01;35:bd=40;33;01:cd=40;33;01:or=40;31;01:mi=00:su=37;41:sg=30;43:ca=30;41:tw=30;42:ow=34;42:st=37;44:ex=01;32:*.tar=01;31:*.tgz=01;31:*.arc=01;31:*.arj=01;31:*.taz=01;31:*.lha=01;31:*.lz4=01;31:*.lzh=01;31:*.lzma=01;31:*.tlz=01;31:*.txz=01;31:*.tzo=01;31:*.t7z=01;31:*.zip=01;31:*.z=01;31:*.Z=01;31:*.dz=01;31:*.gz=01;31:*.lrz=01;31:*.lz=01;31:*.lzo=01;31:*.xz=01;31:*.bz2=01;31:*.bz=01;31:*.tbz=01;31:*.tbz2=01;31:*.tz=01;31:*.deb=01;31:*.rpm=01;31:*.jar=01;31:*.war=01;31:*.ear=01;31:*.sar=01;31:*.rar=01;31:*.alz=01;31:*.ace=01;31:*.zoo=01;31:*.cpio=01;31:*.7z=01;31:*.rz=01;31:*.cab=01;31:*.jpg=01;35:*.jpeg=01;35:*.gif=01;35:*.bmp=01;35:*.pbm=01;35:*.pgm=01;35:*.ppm=01;35:*.tga=01;35:*