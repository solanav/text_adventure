�D            ��    saves/hey.sv    
       Cw@     ����   H�            �    Cw@     ���            ����   ����    ��]a��@���   j@     `���   �D     hey     �D     @���	         save                            hey                             save hey ��]a��`���   R`@     �D     �D      ���   �@     ����   ���           �D     �D     `�,    �q@     �q@     �q@     �q@     �q@     �q@     �q@     �q@     ./log/                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          0q@      ��]a������           0q@     0��            ����   �\"   V@             ����!m`@     ����                   ��]���>m����!m                       �q@     �
    �                    �K     ����   `@      ��]a�����   T@     ����   �D            ��    saves/hey.sv    
       Cw@     ����   H�            �    Cw@     ���            ����   ����    ��]a��@���   j@     `���   �D     hey     �D     @���	         save                            hey                             save hey ��]a��`���   R`@     �D     �D      ���   �@     ����   ���           �D     �D     `�,    �q@     �q@     �q@     �q@     �q@     �q@     �q@     �q@     ./log/                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   P     `@        �$     ��]a�����   x@     ����   �D            ��    saves/hey.sv    
       Cw@     ����   H�            �    Cw@     ���            ����   ����    ��]a��@���   j@     `���   �D     hey     �D     @���	         save                            hey                             save hey ��]a��`���   R`@     �D     �D      ���   �@     ����   ���           �D     �D     `�,    �q@     �q@     �q@     �q@     �q@     �q@     �q@     �q@     ./log/                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          0q@      ��]a������           0q@     0��            ����   �\"   V@             ����!m`@     ����                   ��]���>m����!m                       �q@     �
    �                    `@     ����           �@     ����                 ����   ����           ����   ����   ����     �   '  �   W  �   d  �   n  �   }  �   �  �   �  �   �  �   �  �   �  �   �  �    �   K �   � �   � �   � �    �   > �   r �   � �   � �   � �   ? �   J �   i �   � �   � �   � �   � �      ��     �$     ��]a�����   �@     ����   �D            ��    saves/hey.sv    
       Cw@     ����   H�            �    Cw@     ���            ����   ����    ��]a��@���   j@     `���   �D     hey     �D     @���	         save                            hey                             save hey ��]a��`���   R`@     �D     �D      ���   �@     ����   ���           �D     �D     `�,    �q@     �q@     �q@     �q@     �q@     �q@     �q@     �q@     ./log/                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          0q@      ��]a������           0q@     0��            ����   �\"   V@             ����!m`@     ����                   ��]���>m����!m                       �q@     �
    �                    `@     ����           �@     ����                 ����   ����           ����   ����   ����     �   '  �   W  �   d  �   n  �   }  �   �  �   �  �   �  �   �  �   �  �   �  �    �   K �   � �   � �   � �    �   > �   r �   � �   � �   � �   ? �   J �   i �   � �   � �   � �   � �   
 �    �   3 �   S �   b �   � �      �'     ��]a�����   �@     �p      ��]a��